`define WIDTH		640
`define HEIGHT		480
`define H_FRONT		16
`define H_PULSE		96
`define H_BACK		48
`define V_FRONT		10
`define V_PULSE		2
`define V_BACK		33

`define LINE		`H_PULSE + `H_BACK + `WIDTH + `H_FRONT
`define SCREEN		`V_PULSE + `V_BACK + `HEIGHT + `V_FRONT
